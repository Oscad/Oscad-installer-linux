* eeschema netlist version 1.1 (spice format) creation date: friday 10 january 2014 03:37:10 pm ist

u1  inv nonin vee out vcc port
* The file may be copied, and distributed; however, reselling the 
*  material is illegal

*////////////////////////////////////////////////////////////////////
* For ordering or technical information on these models, contact:
* National Semiconductor's Customer Response Center
*                 7:00 A.M.--7:00 P.M.  U.S. Central Time
*                                (800) 272-9959
* For Applications support, contact the Internet address:
*  amps-apps@galaxy.nsc.com

*//////////////////////////////////////////////////////////
*LM741 OPERATIONAL AMPLIFIER MACRO-MODEL
*//////////////////////////////////////////////////////////
*
* connections:      non-inverting input
*                   |     inverting input
*                   |     |    positive power supply
*                   |     |    |     negative power supply
*                   |     |    |     |    output
*                   |     |    |     |    |
*                   |     |    |     |    |
*                 nonin   inv  vcc  vee  out
*
*Features:
*Improved performance over industry standards
*Plug-in replacement for LM709,LM201,MC1439,748
*Input and output overload protection
*
****************INPUT STAGE**************
*
IOS inv nonin 20N
*^Input offset current
R1 nonin 3 250K
R2 3 inv 250K
I1 4 vee 100U
R3 5 vcc 517
R4 6 vcc 517
Q1 5 inv 4 QX
Q2 6 7 4 QX
*Fp2=2.55 MHz
C4 5 6 60.3614P
*
***********COMMON MODE EFFECT***********
*
I2 vcc vee 1.6MA
*^Quiescent supply current
EOS 7 nonin POLY(1) 16 49 1E-3 1
*Input offset voltage.^
R8 vcc 49 40K
R9 49 vee 40K
*
*********OUTPUT VOLTAGE LIMITING********
V2 vcc 8 1.63
D1 9 8 DX
D2 10 9 DX
V3 10 vee 1.63
*
**************SECOND STAGE**************
*
EH vcc 98 vcc 49 1
G1 98 9 5 6 2.1E-3
*Fp1=5 Hz
R5 98 9 95.493MEG
C3 98 9 333.33P
*
***************POLE STAGE***************
*
*Fp=30 MHz
G3 98 15 9 49 1E-6
R12 98 15 1MEG
C5 98 15 5.3052E-15
*
*********COMMON-MODE ZERO STAGE*********
*
*Fpcm=300 Hz
G4 98 16 3 49 3.1623E-8
L2 98 17 530.5M
R13 17 16 1K
*
**************OUTPUT STAGE**************
*
F6 vee vcc POLY(1) V6 450U 1
E1 vcc 23 vcc 15 1
R16 24 23 25
D5 26 24 DX
V6 26 22 0.65V
R17 23 25 25
D6 25 27 DX
V7 22 27 0.65V
V5 22 21 0.18V
D4 21 15 DX
V4 20 22 0.18V
D3 15 20 DX
L3 22 out 100P
RL3 22 out 100K
*
***************MODELS USED**************
*
.MODEL DX D(IS=1E-15)
.MODEL QX NPN(BF=625)


