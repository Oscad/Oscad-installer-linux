* EESchema Netlist Version 1.1 (Spice format) creation date: Friday 10 January 2014 03:37:10 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
U1  inv nonin VEE out VCC PORT		
U2  inv nonin VEE out VCC opamp1		

.end
